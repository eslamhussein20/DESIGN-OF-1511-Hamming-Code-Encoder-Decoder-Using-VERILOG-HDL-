module HAMMING_ENCODER 
(
input [10:0] ENCODER_IN ,
output [14:0] ENCODER_OUT
);
wire p1 , p2 , p3 , p4 ;
xor (p1,ENCODER_IN[0],ENCODER_IN[1],ENCODER_IN[3],ENCODER_IN[4],ENCODER_IN[6],ENCODER_IN[8],ENCODER_IN[10]);
xor (p2,ENCODER_IN[0],ENCODER_IN[2],ENCODER_IN[3],ENCODER_IN[5],ENCODER_IN[6],ENCODER_IN[9],ENCODER_IN[10]);
xor (p3,ENCODER_IN[1],ENCODER_IN[2],ENCODER_IN[3],ENCODER_IN[7],ENCODER_IN[8],ENCODER_IN[9],ENCODER_IN[10]);
xor (p4,ENCODER_IN[4],ENCODER_IN[5],ENCODER_IN[6],ENCODER_IN[7],ENCODER_IN[8],ENCODER_IN[9],ENCODER_IN[10]);
assign ENCODER_OUT = {ENCODER_IN[10],ENCODER_IN[9] , ENCODER_IN[8],ENCODER_IN[7],ENCODER_IN[6],ENCODER_IN[5],ENCODER_IN[4],p4 , ENCODER_IN[3] , ENCODER_IN[2],ENCODER_IN[1],p3,ENCODER_IN[0],p2,p1 };
endmodule
